`include "defines.vh"

module lsu #(
	parameter XLEN = 32
)(
    input s_load,
    input s_store,
    input funct3
);

endmodule
